library verilog;
use verilog.vl_types.all;
entity tb_CALC1 is
end tb_CALC1;

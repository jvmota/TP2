module CALC1 (
	
);
endmodule

library verilog;
use verilog.vl_types.all;
entity TB_ALU is
end TB_ALU;
